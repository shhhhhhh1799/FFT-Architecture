// `timescale 1ns / 1ps

// 512-point Twiddle Factor ROM 모듈 (<2.7> 형식, signed 9bit 출력)
// addr에 해당하는 twiddle factor를 복소수 형태로 출력함
// 출력은 항상 1클럭 레지스터를 통해 클럭 동기화됨

module twiddle_512 (
    input   clk,
    input [8:0] addr,                 // twiddle 주소 (0~511)
    output signed [8:0] tw_re,       // twiddle의 실수부 (<2.7>)
    output signed [8:0] tw_im        // twiddle의 허수부 (<2.7>)
);

    // 내부 Twiddle Table 정의 (ROM처럼 사용)
    wire [8:0] twf_rom_re[0:511];  // 실수부 테이블
    wire [8:0] twf_rom_im[0:511];  // 허수부 테이블

    // 선택된 twiddle factor
    wire [8:0] mx_re = twf_rom_re[addr];  // MUX로 선택된 실수부
    wire [8:0] mx_im = twf_rom_im[addr];  // MUX로 선택된 허수부

    // 클럭 동기화용 FF
    reg  [8:0] ff_re;         // FF에 저장된 실수부
    reg  [8:0] ff_im;         // FF에 저장된 허수부

    // 클럭 동기화
    always @(posedge clk) begin
        ff_re <= mx_re;
        ff_im <= mx_im;
    end

    // 최종 출력 (무조건 FF 경유)
        assign tw_re = ff_re;
        assign tw_im = ff_im;

    assign  twf_rom_re[  0] = 9'd128;   assign  twf_rom_im[  0] = 0;
    assign  twf_rom_re[  1] = 9'd128;   assign  twf_rom_im[  1] = 0;
    assign  twf_rom_re[  2] = 9'd128;   assign  twf_rom_im[  2] = 0;
    assign  twf_rom_re[  3] = 9'd128;   assign  twf_rom_im[  3] = 0;
    assign  twf_rom_re[  4] = 9'd128;   assign  twf_rom_im[  4] = 0;
    assign  twf_rom_re[  5] = 9'd128;   assign  twf_rom_im[  5] = 0;
    assign  twf_rom_re[  6] = 9'd128;   assign  twf_rom_im[  6] = 0;
    assign  twf_rom_re[  7] = 9'd128;   assign  twf_rom_im[  7] = 0;
    assign  twf_rom_re[  8] = 9'd128;   assign  twf_rom_im[  8] = 0;
    assign  twf_rom_re[  9] = 9'd128;   assign  twf_rom_im[  9] = 0;
    assign  twf_rom_re[ 10] = 9'd128;   assign  twf_rom_im[ 10] = 0;
    assign  twf_rom_re[ 11] = 9'd128;   assign  twf_rom_im[ 11] = 0;
    assign  twf_rom_re[ 12] = 9'd128;   assign  twf_rom_im[ 12] = 0;
    assign  twf_rom_re[ 13] = 9'd128;   assign  twf_rom_im[ 13] = 0;
    assign  twf_rom_re[ 14] = 9'd128;   assign  twf_rom_im[ 14] = 0;
    assign  twf_rom_re[ 15] = 9'd128;   assign  twf_rom_im[ 15] = 0;
    assign  twf_rom_re[ 16] = 9'd128;   assign  twf_rom_im[ 16] = 0;
    assign  twf_rom_re[ 17] = 9'd128;   assign  twf_rom_im[ 17] = 0;
    assign  twf_rom_re[ 18] = 9'd128;   assign  twf_rom_im[ 18] = 0;
    assign  twf_rom_re[ 19] = 9'd128;   assign  twf_rom_im[ 19] = 0;
    assign  twf_rom_re[ 20] = 9'd128;   assign  twf_rom_im[ 20] = 0;
    assign  twf_rom_re[ 21] = 9'd128;   assign  twf_rom_im[ 21] = 0;
    assign  twf_rom_re[ 22] = 9'd128;   assign  twf_rom_im[ 22] = 0;
    assign  twf_rom_re[ 23] = 9'd128;   assign  twf_rom_im[ 23] = 0;
    assign  twf_rom_re[ 24] = 9'd128;   assign  twf_rom_im[ 24] = 0;
    assign  twf_rom_re[ 25] = 9'd128;   assign  twf_rom_im[ 25] = 0;
    assign  twf_rom_re[ 26] = 9'd128;   assign  twf_rom_im[ 26] = 0;
    assign  twf_rom_re[ 27] = 9'd128;   assign  twf_rom_im[ 27] = 0;
    assign  twf_rom_re[ 28] = 9'd128;   assign  twf_rom_im[ 28] = 0;
    assign  twf_rom_re[ 29] = 9'd128;   assign  twf_rom_im[ 29] = 0;
    assign  twf_rom_re[ 30] = 9'd128;   assign  twf_rom_im[ 30] = 0;
    assign  twf_rom_re[ 31] = 9'd128;   assign  twf_rom_im[ 31] = 0;
    assign  twf_rom_re[ 32] = 9'd128;   assign  twf_rom_im[ 32] = 0;
    assign  twf_rom_re[ 33] = 9'd128;   assign  twf_rom_im[ 33] = 0;
    assign  twf_rom_re[ 34] = 9'd128;   assign  twf_rom_im[ 34] = 0;
    assign  twf_rom_re[ 35] = 9'd128;   assign  twf_rom_im[ 35] = 0;
    assign  twf_rom_re[ 36] = 9'd128;   assign  twf_rom_im[ 36] = 0;
    assign  twf_rom_re[ 37] = 9'd128;   assign  twf_rom_im[ 37] = 0;
    assign  twf_rom_re[ 38] = 9'd128;   assign  twf_rom_im[ 38] = 0;
    assign  twf_rom_re[ 39] = 9'd128;   assign  twf_rom_im[ 39] = 0;
    assign  twf_rom_re[ 40] = 9'd128;   assign  twf_rom_im[ 40] = 0;
    assign  twf_rom_re[ 41] = 9'd128;   assign  twf_rom_im[ 41] = 0;
    assign  twf_rom_re[ 42] = 9'd128;   assign  twf_rom_im[ 42] = 0;
    assign  twf_rom_re[ 43] = 9'd128;   assign  twf_rom_im[ 43] = 0;
    assign  twf_rom_re[ 44] = 9'd128;   assign  twf_rom_im[ 44] = 0;
    assign  twf_rom_re[ 45] = 9'd128;   assign  twf_rom_im[ 45] = 0;
    assign  twf_rom_re[ 46] = 9'd128;   assign  twf_rom_im[ 46] = 0;
    assign  twf_rom_re[ 47] = 9'd128;   assign  twf_rom_im[ 47] = 0;
    assign  twf_rom_re[ 48] = 9'd128;   assign  twf_rom_im[ 48] = 0;
    assign  twf_rom_re[ 49] = 9'd128;   assign  twf_rom_im[ 49] = 0;
    assign  twf_rom_re[ 50] = 9'd128;   assign  twf_rom_im[ 50] = 0;
    assign  twf_rom_re[ 51] = 9'd128;   assign  twf_rom_im[ 51] = 0;
    assign  twf_rom_re[ 52] = 9'd128;   assign  twf_rom_im[ 52] = 0;
    assign  twf_rom_re[ 53] = 9'd128;   assign  twf_rom_im[ 53] = 0;
    assign  twf_rom_re[ 54] = 9'd128;   assign  twf_rom_im[ 54] = 0;
    assign  twf_rom_re[ 55] = 9'd128;   assign  twf_rom_im[ 55] = 0;
    assign  twf_rom_re[ 56] = 9'd128;   assign  twf_rom_im[ 56] = 0;
    assign  twf_rom_re[ 57] = 9'd128;   assign  twf_rom_im[ 57] = 0;
    assign  twf_rom_re[ 58] = 9'd128;   assign  twf_rom_im[ 58] = 0;
    assign  twf_rom_re[ 59] = 9'd128;   assign  twf_rom_im[ 59] = 0;
    assign  twf_rom_re[ 60] = 9'd128;   assign  twf_rom_im[ 60] = 0;
    assign  twf_rom_re[ 61] = 9'd128;   assign  twf_rom_im[ 61] = 0;
    assign  twf_rom_re[ 62] = 9'd128;   assign  twf_rom_im[ 62] = 0;
    assign  twf_rom_re[ 63] = 9'd128;   assign  twf_rom_im[ 63] = 0;
    assign  twf_rom_re[ 64] = 9'd128;   assign  twf_rom_im[ 64] = 0;
    assign  twf_rom_re[ 65] = 9'd128;   assign  twf_rom_im[ 65] = -9'd6;
    assign  twf_rom_re[ 66] = 9'd127;   assign  twf_rom_im[ 66] = -9'd13;
    assign  twf_rom_re[ 67] = 9'd127;   assign  twf_rom_im[ 67] = -9'd19;
    assign  twf_rom_re[ 68] = 9'd126;   assign  twf_rom_im[ 68] = -9'd25;
    assign  twf_rom_re[ 69] = 9'd124;   assign  twf_rom_im[ 69] = -9'd31;
    assign  twf_rom_re[ 70] = 9'd122;   assign  twf_rom_im[ 70] = -9'd37;
    assign  twf_rom_re[ 71] = 9'd121;   assign  twf_rom_im[ 71] = -9'd43;
    assign  twf_rom_re[ 72] = 9'd118;   assign  twf_rom_im[ 72] = -9'd49;
    assign  twf_rom_re[ 73] = 9'd116;   assign  twf_rom_im[ 73] = -9'd55;
    assign  twf_rom_re[ 74] = 9'd113;   assign  twf_rom_im[ 74] = -9'd60;
    assign  twf_rom_re[ 75] = 9'd110;   assign  twf_rom_im[ 75] = -9'd66;
    assign  twf_rom_re[ 76] = 9'd106;   assign  twf_rom_im[ 76] = -9'd71;
    assign  twf_rom_re[ 77] = 9'd103;   assign  twf_rom_im[ 77] = -9'd76;
    assign  twf_rom_re[ 78] = 9'd99;    assign  twf_rom_im[ 78] = -9'd81;
    assign  twf_rom_re[ 79] = 9'd95;    assign  twf_rom_im[ 79] = -9'd86;
    assign  twf_rom_re[ 80] = 9'd91;    assign  twf_rom_im[ 80] = -9'd91;
    assign  twf_rom_re[ 81] = 9'd86;    assign  twf_rom_im[ 81] = -9'd95;
    assign  twf_rom_re[ 82] = 9'd81;    assign  twf_rom_im[ 82] = -9'd99;
    assign  twf_rom_re[ 83] = 9'd76;    assign  twf_rom_im[ 83] = -9'd103; 
    assign  twf_rom_re[ 84] = 9'd71;    assign  twf_rom_im[ 84] = -9'd106; 
    assign  twf_rom_re[ 85] = 9'd66;    assign  twf_rom_im[ 85] = -9'd110; 
    assign  twf_rom_re[ 86] = 9'd60;    assign  twf_rom_im[ 86] = -9'd113; 
    assign  twf_rom_re[ 87] = 9'd55;    assign  twf_rom_im[ 87] = -9'd116; 
    assign  twf_rom_re[ 88] = 9'd49;    assign  twf_rom_im[ 88] = -9'd118; 
    assign  twf_rom_re[ 89] = 9'd43;    assign  twf_rom_im[ 89] = -9'd121; 
    assign  twf_rom_re[ 90] = 9'd37;    assign  twf_rom_im[ 90] = -9'd122; 
    assign  twf_rom_re[ 91] = 9'd31;    assign  twf_rom_im[ 91] = -9'd124; 
    assign  twf_rom_re[ 92] = 9'd25;    assign  twf_rom_im[ 92] = -9'd126; 
    assign  twf_rom_re[ 93] = 9'd19;    assign  twf_rom_im[ 93] = -9'd127; 
    assign  twf_rom_re[ 94] = 9'd13;    assign  twf_rom_im[ 94] = -9'd127; 
    assign  twf_rom_re[ 95] = 9'd6;     assign  twf_rom_im[ 95] = -9'd128; 
    assign  twf_rom_re[ 96] = 9'd0;     assign  twf_rom_im[ 96] = -9'd128; 
    assign  twf_rom_re[ 97] = -9'd6;    assign  twf_rom_im[ 97] = -9'd128; 
    assign  twf_rom_re[ 98] = -9'd13;   assign  twf_rom_im[ 98] = -9'd127; 
    assign  twf_rom_re[ 99] = -9'd19;   assign  twf_rom_im[ 99] = -9'd127; 
    assign  twf_rom_re[100] = -9'd25;   assign  twf_rom_im[100] = -9'd126;
    assign  twf_rom_re[101] = -9'd31;   assign  twf_rom_im[101] = -9'd124;
    assign  twf_rom_re[102] = -9'd37;   assign  twf_rom_im[102] = -9'd122;
    assign  twf_rom_re[103] = -9'd43;   assign  twf_rom_im[103] = -9'd121;
    assign  twf_rom_re[104] = -9'd49;   assign  twf_rom_im[104] = -9'd118;
    assign  twf_rom_re[105] = -9'd55;   assign  twf_rom_im[105] = -9'd116;
    assign  twf_rom_re[106] = -9'd60;   assign  twf_rom_im[106] = -9'd113;
    assign  twf_rom_re[107] = -9'd66;   assign  twf_rom_im[107] = -9'd110;
    assign  twf_rom_re[108] = -9'd71;   assign  twf_rom_im[108] = -9'd106;
    assign  twf_rom_re[109] = -9'd76;   assign  twf_rom_im[109] = -9'd103;
    assign  twf_rom_re[110] = -9'd81;   assign  twf_rom_im[110] = -9'd99;
    assign  twf_rom_re[111] = -9'd86;   assign  twf_rom_im[111] = -9'd95;
    assign  twf_rom_re[112] = -9'd91;   assign  twf_rom_im[112] = -9'd91;
    assign  twf_rom_re[113] = -9'd95;   assign  twf_rom_im[113] = -9'd86;
    assign  twf_rom_re[114] = -9'd99;   assign  twf_rom_im[114] = -9'd81;
    assign  twf_rom_re[115] = -9'd103;  assign  twf_rom_im[115] =-9'd76;
    assign  twf_rom_re[116] = -9'd106;  assign  twf_rom_im[116] =-9'd71;
    assign  twf_rom_re[117] = -9'd110;  assign  twf_rom_im[117] =-9'd66;
    assign  twf_rom_re[118] = -9'd113;  assign  twf_rom_im[118] =-9'd60;
    assign  twf_rom_re[119] = -9'd116;  assign  twf_rom_im[119] =-9'd55;
    assign  twf_rom_re[120] = -9'd118;  assign  twf_rom_im[120] =-9'd49;
    assign  twf_rom_re[121] = -9'd121;  assign  twf_rom_im[121] =-9'd43;
    assign  twf_rom_re[122] = -9'd122;  assign  twf_rom_im[122] =-9'd37;
    assign  twf_rom_re[123] = -9'd124;  assign  twf_rom_im[123] =-9'd31;
    assign  twf_rom_re[124] = -9'd126;  assign  twf_rom_im[124] =-9'd25;
    assign  twf_rom_re[125] = -9'd127;  assign  twf_rom_im[125] =-9'd19;
    assign  twf_rom_re[126] = -9'd127;  assign  twf_rom_im[126] =-9'd13;
    assign  twf_rom_re[127] = -9'd128;  assign  twf_rom_im[127] =-9'd6;
    assign  twf_rom_re[128] = 9'd128;   assign  twf_rom_im[128] = 0;
    assign  twf_rom_re[129] = 9'd128;   assign  twf_rom_im[129] = -9'd3;
    assign  twf_rom_re[130] = 9'd128;   assign  twf_rom_im[130] = -9'd6;
    assign  twf_rom_re[131] = 9'd128;   assign  twf_rom_im[131] = -9'd9;
    assign  twf_rom_re[132] = 9'd127;   assign  twf_rom_im[132] = -9'd13;
    assign  twf_rom_re[133] = 9'd127;   assign  twf_rom_im[133] = -9'd16;
    assign  twf_rom_re[134] = 9'd127;   assign  twf_rom_im[134] = -9'd19;
    assign  twf_rom_re[135] = 9'd126;   assign  twf_rom_im[135] = -9'd22;
    assign  twf_rom_re[136] = 9'd126;   assign  twf_rom_im[136] = -9'd25;
    assign  twf_rom_re[137] = 9'd125;   assign  twf_rom_im[137] = -9'd28;
    assign  twf_rom_re[138] = 9'd124;   assign  twf_rom_im[138] = -9'd31;
    assign  twf_rom_re[139] = 9'd123;   assign  twf_rom_im[139] = -9'd34;
    assign  twf_rom_re[140] = 9'd122;   assign  twf_rom_im[140] = -9'd37;
    assign  twf_rom_re[141] = 9'd122;   assign  twf_rom_im[141] = -9'd40;
    assign  twf_rom_re[142] = 9'd121;   assign  twf_rom_im[142] = -9'd43;
    assign  twf_rom_re[143] = 9'd119;   assign  twf_rom_im[143] = -9'd46;
    assign  twf_rom_re[144] = 9'd118;   assign  twf_rom_im[144] = -9'd49;
    assign  twf_rom_re[145] = 9'd117;   assign  twf_rom_im[145] = -9'd52;
    assign  twf_rom_re[146] = 9'd116;   assign  twf_rom_im[146] = -9'd55;
    assign  twf_rom_re[147] = 9'd114;   assign  twf_rom_im[147] = -9'd58;
    assign  twf_rom_re[148] = 9'd113;   assign  twf_rom_im[148] = -9'd60;
    assign  twf_rom_re[149] = 9'd111;   assign  twf_rom_im[149] = -9'd63;
    assign  twf_rom_re[150] = 9'd110;   assign  twf_rom_im[150] = -9'd66;
    assign  twf_rom_re[151] = 9'd108;   assign  twf_rom_im[151] = -9'd68;
    assign  twf_rom_re[152] = 9'd106;   assign  twf_rom_im[152] = -9'd71;
    assign  twf_rom_re[153] = 9'd105;   assign  twf_rom_im[153] = -9'd74;
    assign  twf_rom_re[154] = 9'd103;   assign  twf_rom_im[154] = -9'd76;
    assign  twf_rom_re[155] = 9'd101;   assign  twf_rom_im[155] = -9'd79;
    assign  twf_rom_re[156] = 9'd99;    assign  twf_rom_im[156] = -9'd81;
    assign  twf_rom_re[157] = 9'd97;    assign  twf_rom_im[157] = -9'd84;
    assign  twf_rom_re[158] = 9'd95;    assign  twf_rom_im[158] = -9'd86;
    assign  twf_rom_re[159] = 9'd93;    assign  twf_rom_im[159] = -9'd88;
    assign  twf_rom_re[160] = 9'd91;    assign  twf_rom_im[160] = -9'd91;
    assign  twf_rom_re[161] = 9'd88;    assign  twf_rom_im[161] = -9'd93;
    assign  twf_rom_re[162] = 9'd86;    assign  twf_rom_im[162] = -9'd95;
    assign  twf_rom_re[163] = 9'd84;    assign  twf_rom_im[163] = -9'd97;
    assign  twf_rom_re[164] = 9'd81;    assign  twf_rom_im[164] = -9'd99;
    assign  twf_rom_re[165] = 9'd79;    assign  twf_rom_im[165] = -9'd101;
    assign  twf_rom_re[166] = 9'd76;    assign  twf_rom_im[166] = -9'd103;
    assign  twf_rom_re[167] = 9'd74;    assign  twf_rom_im[167] = -9'd105;
    assign  twf_rom_re[168] = 9'd71;    assign  twf_rom_im[168] = -9'd106;
    assign  twf_rom_re[169] = 9'd68;    assign  twf_rom_im[169] = -9'd108;
    assign  twf_rom_re[170] = 9'd66;    assign  twf_rom_im[170] = -9'd110;
    assign  twf_rom_re[171] = 9'd63;    assign  twf_rom_im[171] = -9'd111;
    assign  twf_rom_re[172] = 9'd60;    assign  twf_rom_im[172] = -9'd113;
    assign  twf_rom_re[173] = 9'd58;    assign  twf_rom_im[173] = -9'd114;
    assign  twf_rom_re[174] = 9'd55;    assign  twf_rom_im[174] = -9'd116;
    assign  twf_rom_re[175] = 9'd52;    assign  twf_rom_im[175] = -9'd117;
    assign  twf_rom_re[176] = 9'd49;    assign  twf_rom_im[176] = -9'd118;
    assign  twf_rom_re[177] = 9'd46;    assign  twf_rom_im[177] = -9'd119;
    assign  twf_rom_re[178] = 9'd43;    assign  twf_rom_im[178] = -9'd121;
    assign  twf_rom_re[179] = 9'd40;    assign  twf_rom_im[179] = -9'd122;
    assign  twf_rom_re[180] = 9'd37;    assign  twf_rom_im[180] = -9'd122;
    assign  twf_rom_re[181] = 9'd34;    assign  twf_rom_im[181] = -9'd123;
    assign  twf_rom_re[182] = 9'd31;    assign  twf_rom_im[182] = -9'd124;
    assign  twf_rom_re[183] = 9'd28;    assign  twf_rom_im[183] = -9'd125;
    assign  twf_rom_re[184] = 9'd25;    assign  twf_rom_im[184] = -9'd126;
    assign  twf_rom_re[185] = 9'd22;    assign  twf_rom_im[185] = -9'd126;
    assign  twf_rom_re[186] = 9'd19;    assign  twf_rom_im[186] = -9'd127;
    assign  twf_rom_re[187] = 9'd16;    assign  twf_rom_im[187] = -9'd127;
    assign  twf_rom_re[188] = 9'd13;    assign  twf_rom_im[188] = -9'd127;
    assign  twf_rom_re[189] = 9'd9;     assign  twf_rom_im[189] = -9'd128;
    assign  twf_rom_re[190] = 9'd6;     assign  twf_rom_im[190] = -9'd128;
    assign  twf_rom_re[191] = 9'd3;     assign  twf_rom_im[191] = -9'd128;
    assign  twf_rom_re[192] = 9'd128;   assign  twf_rom_im[192] = 0;
    assign  twf_rom_re[193] = 9'd128;   assign  twf_rom_im[193] = -9'd9;
    assign  twf_rom_re[194] = 9'd127;   assign  twf_rom_im[194] = -9'd19;
    assign  twf_rom_re[195] = 9'd125;   assign  twf_rom_im[195] = -9'd28;
    assign  twf_rom_re[196] = 9'd122;   assign  twf_rom_im[196] = -9'd37;
    assign  twf_rom_re[197] = 9'd119;   assign  twf_rom_im[197] = -9'd46;
    assign  twf_rom_re[198] = 9'd116;   assign  twf_rom_im[198] = -9'd55;
    assign  twf_rom_re[199] = 9'd111;   assign  twf_rom_im[199] = -9'd63;
    assign  twf_rom_re[200] = 9'd106;   assign  twf_rom_im[200] = -9'd71;
    assign  twf_rom_re[201] = 9'd101;   assign  twf_rom_im[201] = -9'd79;
    assign  twf_rom_re[202] = 9'd95;    assign  twf_rom_im[202] = -9'd86;
    assign  twf_rom_re[203] = 9'd88;    assign  twf_rom_im[203] = -9'd93;
    assign  twf_rom_re[204] = 9'd81;    assign  twf_rom_im[204] = -9'd99;
    assign  twf_rom_re[205] = 9'd74;    assign  twf_rom_im[205] = -9'd105;
    assign  twf_rom_re[206] = 9'd66;    assign  twf_rom_im[206] = -9'd110;
    assign  twf_rom_re[207] = 9'd58;    assign  twf_rom_im[207] = -9'd114;
    assign  twf_rom_re[208] = 9'd49;    assign  twf_rom_im[208] = -9'd118;
    assign  twf_rom_re[209] = 9'd40;    assign  twf_rom_im[209] = -9'd122;
    assign  twf_rom_re[210] = 9'd31;    assign  twf_rom_im[210] = -9'd124;
    assign  twf_rom_re[211] = 9'd22;    assign  twf_rom_im[211] = -9'd126;
    assign  twf_rom_re[212] = 9'd13;    assign  twf_rom_im[212] = -9'd127;
    assign  twf_rom_re[213] = 9'd3;     assign  twf_rom_im[213] = -9'd128;
    assign  twf_rom_re[214] = -9'd6;    assign  twf_rom_im[214] = -9'd128;
    assign  twf_rom_re[215] = -9'd16;   assign  twf_rom_im[215] = -9'd127;
    assign  twf_rom_re[216] = -9'd25;   assign  twf_rom_im[216] = -9'd126;
    assign  twf_rom_re[217] = -9'd34;   assign  twf_rom_im[217] = -9'd123;
    assign  twf_rom_re[218] = -9'd43;   assign  twf_rom_im[218] = -9'd121;
    assign  twf_rom_re[219] = -9'd52;   assign  twf_rom_im[219] = -9'd117;
    assign  twf_rom_re[220] = -9'd60;   assign  twf_rom_im[220] = -9'd113;
    assign  twf_rom_re[221] = -9'd68;   assign  twf_rom_im[221] = -9'd108;
    assign  twf_rom_re[222] = -9'd76;   assign  twf_rom_im[222] = -9'd103;
    assign  twf_rom_re[223] = -9'd84;   assign  twf_rom_im[223] = -9'd97;
    assign  twf_rom_re[224] = -9'd91;   assign  twf_rom_im[224] = -9'd91;
    assign  twf_rom_re[225] = -9'd97;   assign  twf_rom_im[225] = -9'd84;
    assign  twf_rom_re[226] = -9'd103;  assign  twf_rom_im[226] = -9'd76;
    assign  twf_rom_re[227] = -9'd108;  assign  twf_rom_im[227] = -9'd68;
    assign  twf_rom_re[228] = -9'd113;  assign  twf_rom_im[228] = -9'd60;
    assign  twf_rom_re[229] = -9'd117;  assign  twf_rom_im[229] = -9'd52;
    assign  twf_rom_re[230] = -9'd121;  assign  twf_rom_im[230] = -9'd43;
    assign  twf_rom_re[231] = -9'd123;  assign  twf_rom_im[231] = -9'd34;
    assign  twf_rom_re[232] = -9'd126;  assign  twf_rom_im[232] = -9'd25;
    assign  twf_rom_re[233] = -9'd127;  assign  twf_rom_im[233] = -9'd16;
    assign  twf_rom_re[234] = -9'd128;  assign  twf_rom_im[234] = -9'd6;
    assign  twf_rom_re[235] = -9'd128;  assign  twf_rom_im[235] = 9'd3;
    assign  twf_rom_re[236] = -9'd127;  assign  twf_rom_im[236] = 9'd13;
    assign  twf_rom_re[237] = -9'd126;  assign  twf_rom_im[237] = 9'd22;
    assign  twf_rom_re[238] = -9'd124;  assign  twf_rom_im[238] = 9'd31;
    assign  twf_rom_re[239] = -9'd122;  assign  twf_rom_im[239] = 9'd40;
    assign  twf_rom_re[240] = -9'd118;  assign  twf_rom_im[240] = 9'd49;
    assign  twf_rom_re[241] = -9'd114;  assign  twf_rom_im[241] = 9'd58;
    assign  twf_rom_re[242] = -9'd110;  assign  twf_rom_im[242] = 9'd66;
    assign  twf_rom_re[243] = -9'd105;  assign  twf_rom_im[243] = 9'd74;
    assign  twf_rom_re[244] = -9'd99;   assign  twf_rom_im[244] = 9'd81;
    assign  twf_rom_re[245] = -9'd93;   assign  twf_rom_im[245] = 9'd88;
    assign  twf_rom_re[246] = -9'd86;   assign  twf_rom_im[246] = 9'd95;
    assign  twf_rom_re[247] = -9'd79;   assign  twf_rom_im[247] = 9'd101;
    assign  twf_rom_re[248] = -9'd71;   assign  twf_rom_im[248] = 9'd106;
    assign  twf_rom_re[249] = -9'd63;   assign  twf_rom_im[249] = 9'd111;
    assign  twf_rom_re[250] = -9'd55;   assign  twf_rom_im[250] = 9'd116;
    assign  twf_rom_re[251] = -9'd46;   assign  twf_rom_im[251] = 9'd119;
    assign  twf_rom_re[252] = -9'd37;   assign  twf_rom_im[252] = 9'd122;
    assign  twf_rom_re[253] = -9'd28;   assign  twf_rom_im[253] = 9'd125;
    assign  twf_rom_re[254] = -9'd19;   assign  twf_rom_im[254] = 9'd127;
    assign  twf_rom_re[255] = -9'd9;    assign  twf_rom_im[255] = 9'd128;
    assign  twf_rom_re[256] = 9'd128;   assign  twf_rom_im[256] = 0;
    assign  twf_rom_re[257] = 9'd128;   assign  twf_rom_im[257] = -9'd2;
    assign  twf_rom_re[258] = 9'd128;   assign  twf_rom_im[258] = -9'd3;
    assign  twf_rom_re[259] = 9'd128;   assign  twf_rom_im[259] = -9'd5;
    assign  twf_rom_re[260] = 9'd128;   assign  twf_rom_im[260] = -9'd6;
    assign  twf_rom_re[261] = 9'd128;   assign  twf_rom_im[261] = -9'd8;
    assign  twf_rom_re[262] = 9'd128;   assign  twf_rom_im[262] = -9'd9;
    assign  twf_rom_re[263] = 9'd128;   assign  twf_rom_im[263] = -9'd11;
    assign  twf_rom_re[264] = 9'd127;   assign  twf_rom_im[264] = -9'd13;
    assign  twf_rom_re[265] = 9'd127;   assign  twf_rom_im[265] = -9'd14;
    assign  twf_rom_re[266] = 9'd127;   assign  twf_rom_im[266] = -9'd16;
    assign  twf_rom_re[267] = 9'd127;   assign  twf_rom_im[267] = -9'd17;
    assign  twf_rom_re[268] = 9'd127;   assign  twf_rom_im[268] = -9'd19;
    assign  twf_rom_re[269] = 9'd126;   assign  twf_rom_im[269] = -9'd20;
    assign  twf_rom_re[270] = 9'd126;   assign  twf_rom_im[270] = -9'd22;
    assign  twf_rom_re[271] = 9'd126;   assign  twf_rom_im[271] = -9'd23;
    assign  twf_rom_re[272] = 9'd126;   assign  twf_rom_im[272] = -9'd25;
    assign  twf_rom_re[273] = 9'd125;   assign  twf_rom_im[273] = -9'd27;
    assign  twf_rom_re[274] = 9'd125;   assign  twf_rom_im[274] = -9'd28;
    assign  twf_rom_re[275] = 9'd125;   assign  twf_rom_im[275] = -9'd30;
    assign  twf_rom_re[276] = 9'd124;   assign  twf_rom_im[276] = -9'd31;
    assign  twf_rom_re[277] = 9'd124;   assign  twf_rom_im[277] = -9'd33;
    assign  twf_rom_re[278] = 9'd123;   assign  twf_rom_im[278] = -9'd34;
    assign  twf_rom_re[279] = 9'd123;   assign  twf_rom_im[279] = -9'd36;
    assign  twf_rom_re[280] = 9'd122;   assign  twf_rom_im[280] = -9'd37;
    assign  twf_rom_re[281] = 9'd122;   assign  twf_rom_im[281] = -9'd39;
    assign  twf_rom_re[282] = 9'd122;   assign  twf_rom_im[282] = -9'd40;
    assign  twf_rom_re[283] = 9'd121;   assign  twf_rom_im[283] = -9'd42;
    assign  twf_rom_re[284] = 9'd121;   assign  twf_rom_im[284] = -9'd43;
    assign  twf_rom_re[285] = 9'd120;   assign  twf_rom_im[285] = -9'd45;
    assign  twf_rom_re[286] = 9'd119;   assign  twf_rom_im[286] = -9'd46;
    assign  twf_rom_re[287] = 9'd119;   assign  twf_rom_im[287] = -9'd48;
    assign  twf_rom_re[288] = 9'd118;   assign  twf_rom_im[288] = -9'd49;
    assign  twf_rom_re[289] = 9'd118;   assign  twf_rom_im[289] = -9'd50;
    assign  twf_rom_re[290] = 9'd117;   assign  twf_rom_im[290] = -9'd52;
    assign  twf_rom_re[291] = 9'd116;   assign  twf_rom_im[291] = -9'd53;
    assign  twf_rom_re[292] = 9'd116;   assign  twf_rom_im[292] = -9'd55;
    assign  twf_rom_re[293] = 9'd115;   assign  twf_rom_im[293] = -9'd56;
    assign  twf_rom_re[294] = 9'd114;   assign  twf_rom_im[294] = -9'd58;
    assign  twf_rom_re[295] = 9'd114;   assign  twf_rom_im[295] = -9'd59;
    assign  twf_rom_re[296] = 9'd113;   assign  twf_rom_im[296] = -9'd60;
    assign  twf_rom_re[297] = 9'd112;   assign  twf_rom_im[297] = -9'd62;
    assign  twf_rom_re[298] = 9'd111;   assign  twf_rom_im[298] = -9'd63;
    assign  twf_rom_re[299] = 9'd111;   assign  twf_rom_im[299] = -9'd64;
    assign  twf_rom_re[300] = 9'd110;   assign  twf_rom_im[300] = -9'd66;
    assign  twf_rom_re[301] = 9'd109;   assign  twf_rom_im[301] = -9'd67;
    assign  twf_rom_re[302] = 9'd108;   assign  twf_rom_im[302] = -9'd68;
    assign  twf_rom_re[303] = 9'd107;   assign  twf_rom_im[303] = -9'd70;
    assign  twf_rom_re[304] = 9'd106;   assign  twf_rom_im[304] = -9'd71;
    assign  twf_rom_re[305] = 9'd106;   assign  twf_rom_im[305] = -9'd72;
    assign  twf_rom_re[306] = 9'd105;   assign  twf_rom_im[306] = -9'd74;
    assign  twf_rom_re[307] = 9'd104;   assign  twf_rom_im[307] = -9'd75;
    assign  twf_rom_re[308] = 9'd103;   assign  twf_rom_im[308] = -9'd76;
    assign  twf_rom_re[309] = 9'd102;   assign  twf_rom_im[309] = -9'd78;
    assign  twf_rom_re[310] = 9'd101;   assign  twf_rom_im[310] = -9'd79;
    assign  twf_rom_re[311] = 9'd100;   assign  twf_rom_im[311] = -9'd80;
    assign  twf_rom_re[312] = 9'd99;    assign  twf_rom_im[312] = -9'd81;
    assign  twf_rom_re[313] = 9'd98;    assign  twf_rom_im[313] = -9'd82;
    assign  twf_rom_re[314] = 9'd97;    assign  twf_rom_im[314] = -9'd84;
    assign  twf_rom_re[315] = 9'd96;    assign  twf_rom_im[315] = -9'd85;
    assign  twf_rom_re[316] = 9'd95;    assign  twf_rom_im[316] = -9'd86;
    assign  twf_rom_re[317] = 9'd94;    assign  twf_rom_im[317] = -9'd87;
    assign  twf_rom_re[318] = 9'd93;    assign  twf_rom_im[318] = -9'd88;
    assign  twf_rom_re[319] = 9'd92;    assign  twf_rom_im[319] = -9'd89;
    assign  twf_rom_re[320] = 9'd128;   assign  twf_rom_im[320] = 0;
    assign  twf_rom_re[321] = 9'd128;   assign  twf_rom_im[321] = -9'd8;
    assign  twf_rom_re[322] = 9'd127;   assign  twf_rom_im[322] = -9'd16;
    assign  twf_rom_re[323] = 9'd126;   assign  twf_rom_im[323] = -9'd23;
    assign  twf_rom_re[324] = 9'd124;   assign  twf_rom_im[324] = -9'd31;
    assign  twf_rom_re[325] = 9'd122;   assign  twf_rom_im[325] = -9'd39;
    assign  twf_rom_re[326] = 9'd119;   assign  twf_rom_im[326] = -9'd46;
    assign  twf_rom_re[327] = 9'd116;   assign  twf_rom_im[327] = -9'd53;
    assign  twf_rom_re[328] = 9'd113;   assign  twf_rom_im[328] = -9'd60;
    assign  twf_rom_re[329] = 9'd109;   assign  twf_rom_im[329] = -9'd67;
    assign  twf_rom_re[330] = 9'd105;   assign  twf_rom_im[330] = -9'd74;
    assign  twf_rom_re[331] = 9'd100;   assign  twf_rom_im[331] = -9'd80;
    assign  twf_rom_re[332] = 9'd95;    assign  twf_rom_im[332] = -9'd86;
    assign  twf_rom_re[333] = 9'd89;    assign  twf_rom_im[333] = -9'd92;
    assign  twf_rom_re[334] = 9'd84;    assign  twf_rom_im[334] = -9'd97;
    assign  twf_rom_re[335] = 9'd78;    assign  twf_rom_im[335] = -9'd102;
    assign  twf_rom_re[336] = 9'd71;    assign  twf_rom_im[336] = -9'd106;
    assign  twf_rom_re[337] = 9'd64;    assign  twf_rom_im[337] = -9'd111;
    assign  twf_rom_re[338] = 9'd58;    assign  twf_rom_im[338] = -9'd114;
    assign  twf_rom_re[339] = 9'd50;    assign  twf_rom_im[339] = -9'd118;
    assign  twf_rom_re[340] = 9'd43;    assign  twf_rom_im[340] = -9'd121;
    assign  twf_rom_re[341] = 9'd36;    assign  twf_rom_im[341] = -9'd123;
    assign  twf_rom_re[342] = 9'd28;    assign  twf_rom_im[342] = -9'd125;
    assign  twf_rom_re[343] = 9'd20;    assign  twf_rom_im[343] = -9'd126;
    assign  twf_rom_re[344] = 9'd13;    assign  twf_rom_im[344] = -9'd127;
    assign  twf_rom_re[345] = 9'd5;     assign  twf_rom_im[345] = -9'd128;
    assign  twf_rom_re[346] = -9'd3;    assign  twf_rom_im[346] = -9'd128;
    assign  twf_rom_re[347] = -9'd11;   assign  twf_rom_im[347] = -9'd128;
    assign  twf_rom_re[348] = -9'd19;   assign  twf_rom_im[348] = -9'd127;
    assign  twf_rom_re[349] = -9'd27;   assign  twf_rom_im[349] = -9'd125;
    assign  twf_rom_re[350] = -9'd34;   assign  twf_rom_im[350] = -9'd123;
    assign  twf_rom_re[351] = -9'd42;   assign  twf_rom_im[351] = -9'd121;
    assign  twf_rom_re[352] = -9'd49;   assign  twf_rom_im[352] = -9'd118;
    assign  twf_rom_re[353] = -9'd56;   assign  twf_rom_im[353] = -9'd115;
    assign  twf_rom_re[354] = -9'd63;   assign  twf_rom_im[354] = -9'd111;
    assign  twf_rom_re[355] = -9'd70;   assign  twf_rom_im[355] = -9'd107;
    assign  twf_rom_re[356] = -9'd76;   assign  twf_rom_im[356] = -9'd103;
    assign  twf_rom_re[357] = -9'd82;   assign  twf_rom_im[357] = -9'd98;
    assign  twf_rom_re[358] = -9'd88;   assign  twf_rom_im[358] = -9'd93;
    assign  twf_rom_re[359] = -9'd94;   assign  twf_rom_im[359] = -9'd87;
    assign  twf_rom_re[360] = -9'd99;   assign  twf_rom_im[360] = -9'd81;
    assign  twf_rom_re[361] = -9'd104;  assign  twf_rom_im[361] = -9'd75;
    assign  twf_rom_re[362] = -9'd108;  assign  twf_rom_im[362] = -9'd68;
    assign  twf_rom_re[363] = -9'd112;  assign  twf_rom_im[363] = -9'd62;
    assign  twf_rom_re[364] = -9'd116;  assign  twf_rom_im[364] = -9'd55;
    assign  twf_rom_re[365] = -9'd119;  assign  twf_rom_im[365] = -9'd48;
    assign  twf_rom_re[366] = -9'd122;  assign  twf_rom_im[366] = -9'd40;
    assign  twf_rom_re[367] = -9'd124;  assign  twf_rom_im[367] = -9'd33;
    assign  twf_rom_re[368] = -9'd126;  assign  twf_rom_im[368] = -9'd25;
    assign  twf_rom_re[369] = -9'd127;  assign  twf_rom_im[369] = -9'd17;
    assign  twf_rom_re[370] = -9'd128;  assign  twf_rom_im[370] = -9'd9;
    assign  twf_rom_re[371] = -9'd128;  assign  twf_rom_im[371] = -9'd2;
    assign  twf_rom_re[372] = -9'd128;  assign  twf_rom_im[372] = 9'd6;
    assign  twf_rom_re[373] = -9'd127;  assign  twf_rom_im[373] = 9'd14;
    assign  twf_rom_re[374] = -9'd126;  assign  twf_rom_im[374] = 9'd22;
    assign  twf_rom_re[375] = -9'd125;  assign  twf_rom_im[375] = 9'd30;
    assign  twf_rom_re[376] = -9'd122;  assign  twf_rom_im[376] = 9'd37;
    assign  twf_rom_re[377] = -9'd120;  assign  twf_rom_im[377] = 9'd45;
    assign  twf_rom_re[378] = -9'd117;  assign  twf_rom_im[378] = 9'd52;
    assign  twf_rom_re[379] = -9'd114;  assign  twf_rom_im[379] = 9'd59;
    assign  twf_rom_re[380] = -9'd110;  assign  twf_rom_im[380] = 9'd66;
    assign  twf_rom_re[381] = -9'd106;  assign  twf_rom_im[381] = 9'd72;
    assign  twf_rom_re[382] = -9'd101;  assign  twf_rom_im[382] = 9'd79;
    assign  twf_rom_re[383] = -9'd96;   assign  twf_rom_im[383] = 9'd85;
    assign  twf_rom_re[384] = 9'd128;   assign  twf_rom_im[384] = 9'd0;
    assign  twf_rom_re[385] = 9'd128;   assign  twf_rom_im[385] = -9'd5;
    assign  twf_rom_re[386] = 9'd128;   assign  twf_rom_im[386] = -9'd9;
    assign  twf_rom_re[387] = 9'd127;   assign  twf_rom_im[387] = -9'd14;
    assign  twf_rom_re[388] = 9'd127;   assign  twf_rom_im[388] = -9'd19;
    assign  twf_rom_re[389] = 9'd126;   assign  twf_rom_im[389] = -9'd23;
    assign  twf_rom_re[390] = 9'd125;   assign  twf_rom_im[390] = -9'd28;
    assign  twf_rom_re[391] = 9'd124;   assign  twf_rom_im[391] = -9'd33;
    assign  twf_rom_re[392] = 9'd122;   assign  twf_rom_im[392] = -9'd37;
    assign  twf_rom_re[393] = 9'd121;   assign  twf_rom_im[393] = -9'd42;
    assign  twf_rom_re[394] = 9'd119;   assign  twf_rom_im[394] = -9'd46;
    assign  twf_rom_re[395] = 9'd118;   assign  twf_rom_im[395] = -9'd50;
    assign  twf_rom_re[396] = 9'd116;   assign  twf_rom_im[396] = -9'd55;
    assign  twf_rom_re[397] = 9'd114;   assign  twf_rom_im[397] = -9'd59;
    assign  twf_rom_re[398] = 9'd111;   assign  twf_rom_im[398] = -9'd63;
    assign  twf_rom_re[399] = 9'd109;   assign  twf_rom_im[399] = -9'd67;
    assign  twf_rom_re[400] = 9'd106;   assign  twf_rom_im[400] = -9'd71;
    assign  twf_rom_re[401] = 9'd104;   assign  twf_rom_im[401] = -9'd75;
    assign  twf_rom_re[402] = 9'd101;   assign  twf_rom_im[402] = -9'd79;
    assign  twf_rom_re[403] = 9'd98;    assign  twf_rom_im[403] = -9'd82;
    assign  twf_rom_re[404] = 9'd95;    assign  twf_rom_im[404] = -9'd86;
    assign  twf_rom_re[405] = 9'd92;    assign  twf_rom_im[405] = -9'd89;
    assign  twf_rom_re[406] = 9'd88;    assign  twf_rom_im[406] = -9'd93;
    assign  twf_rom_re[407] = 9'd85;    assign  twf_rom_im[407] = -9'd96;
    assign  twf_rom_re[408] = 9'd81;    assign  twf_rom_im[408] = -9'd99;
    assign  twf_rom_re[409] = 9'd78;    assign  twf_rom_im[409] = -9'd102;
    assign  twf_rom_re[410] = 9'd74;    assign  twf_rom_im[410] = -9'd105;
    assign  twf_rom_re[411] = 9'd70;    assign  twf_rom_im[411] = -9'd107;
    assign  twf_rom_re[412] = 9'd66;    assign  twf_rom_im[412] = -9'd110;
    assign  twf_rom_re[413] = 9'd62;    assign  twf_rom_im[413] = -9'd112;
    assign  twf_rom_re[414] = 9'd58;    assign  twf_rom_im[414] = -9'd114;
    assign  twf_rom_re[415] = 9'd53;    assign  twf_rom_im[415] = -9'd116;
    assign  twf_rom_re[416] = 9'd49;    assign  twf_rom_im[416] = -9'd118;
    assign  twf_rom_re[417] = 9'd45;    assign  twf_rom_im[417] = -9'd120;
    assign  twf_rom_re[418] = 9'd40;    assign  twf_rom_im[418] = -9'd122;
    assign  twf_rom_re[419] = 9'd36;    assign  twf_rom_im[419] = -9'd123;
    assign  twf_rom_re[420] = 9'd31;    assign  twf_rom_im[420] = -9'd124;
    assign  twf_rom_re[421] = 9'd27;    assign  twf_rom_im[421] = -9'd125;
    assign  twf_rom_re[422] = 9'd22;    assign  twf_rom_im[422] = -9'd126;
    assign  twf_rom_re[423] = 9'd17;    assign  twf_rom_im[423] = -9'd127;
    assign  twf_rom_re[424] = 9'd13;    assign  twf_rom_im[424] = -9'd127;
    assign  twf_rom_re[425] = 9'd8;     assign  twf_rom_im[425] = -9'd128;
    assign  twf_rom_re[426] = 9'd3;     assign  twf_rom_im[426] = -9'd128;
    assign  twf_rom_re[427] = -9'd2;    assign  twf_rom_im[427] = -9'd128;
    assign  twf_rom_re[428] = -9'd6;    assign  twf_rom_im[428] = -9'd128;
    assign  twf_rom_re[429] = -9'd11;   assign  twf_rom_im[429] = -9'd128;
    assign  twf_rom_re[430] = -9'd16;   assign  twf_rom_im[430] = -9'd127;
    assign  twf_rom_re[431] = -9'd20;   assign  twf_rom_im[431] = -9'd126;
    assign  twf_rom_re[432] = -9'd25;   assign  twf_rom_im[432] = -9'd126;
    assign  twf_rom_re[433] = -9'd30;   assign  twf_rom_im[433] = -9'd125;
    assign  twf_rom_re[434] = -9'd34;   assign  twf_rom_im[434] = -9'd123;
    assign  twf_rom_re[435] = -9'd39;   assign  twf_rom_im[435] = -9'd122;
    assign  twf_rom_re[436] = -9'd43;   assign  twf_rom_im[436] = -9'd121;
    assign  twf_rom_re[437] = -9'd48;   assign  twf_rom_im[437] = -9'd119;
    assign  twf_rom_re[438] = -9'd52;   assign  twf_rom_im[438] = -9'd117;
    assign  twf_rom_re[439] = -9'd56;   assign  twf_rom_im[439] = -9'd115;
    assign  twf_rom_re[440] = -9'd60;   assign  twf_rom_im[440] = -9'd113;
    assign  twf_rom_re[441] = -9'd64;   assign  twf_rom_im[441] = -9'd111;
    assign  twf_rom_re[442] = -9'd68;   assign  twf_rom_im[442] = -9'd108;
    assign  twf_rom_re[443] = -9'd72;   assign  twf_rom_im[443] = -9'd106;
    assign  twf_rom_re[444] = -9'd76;   assign  twf_rom_im[444] = -9'd103;
    assign  twf_rom_re[445] = -9'd80;   assign  twf_rom_im[445] = -9'd100;
    assign  twf_rom_re[446] = -9'd84;   assign  twf_rom_im[446] = -9'd97;
    assign  twf_rom_re[447] = -9'd87;   assign  twf_rom_im[447] = -9'd94;
    assign  twf_rom_re[448] = 9'd128;   assign  twf_rom_im[448] = 0;
    assign  twf_rom_re[449] = 9'd128;   assign  twf_rom_im[449] = -9'd11;
    assign  twf_rom_re[450] = 9'd126;   assign  twf_rom_im[450] = -9'd22;
    assign  twf_rom_re[451] = 9'd124;   assign  twf_rom_im[451] = -9'd33;
    assign  twf_rom_re[452] = 9'd121;   assign  twf_rom_im[452] = -9'd43;
    assign  twf_rom_re[453] = 9'd116;   assign  twf_rom_im[453] = -9'd53;
    assign  twf_rom_re[454] = 9'd111;   assign  twf_rom_im[454] = -9'd63;
    assign  twf_rom_re[455] = 9'd106;   assign  twf_rom_im[455] = -9'd72;
    assign  twf_rom_re[456] = 9'd99;    assign  twf_rom_im[456] = -9'd81;
    assign  twf_rom_re[457] = 9'd92;    assign  twf_rom_im[457] = -9'd89;
    assign  twf_rom_re[458] = 9'd84;    assign  twf_rom_im[458] = -9'd97;
    assign  twf_rom_re[459] = 9'd75;    assign  twf_rom_im[459] = -9'd104;
    assign  twf_rom_re[460] = 9'd66;    assign  twf_rom_im[460] = -9'd110;
    assign  twf_rom_re[461] = 9'd56;    assign  twf_rom_im[461] = -9'd115;
    assign  twf_rom_re[462] = 9'd46;    assign  twf_rom_im[462] = -9'd119;
    assign  twf_rom_re[463] = 9'd36;    assign  twf_rom_im[463] = -9'd123;
    assign  twf_rom_re[464] = 9'd25;    assign  twf_rom_im[464] = -9'd126;
    assign  twf_rom_re[465] = 9'd14;    assign  twf_rom_im[465] = -9'd127;
    assign  twf_rom_re[466] = 9'd3;     assign  twf_rom_im[466] = -9'd128;
    assign  twf_rom_re[467] = -9'd8;    assign  twf_rom_im[467] = -9'd128;
    assign  twf_rom_re[468] = -9'd19;   assign  twf_rom_im[468] = -9'd127;
    assign  twf_rom_re[469] = -9'd30;   assign  twf_rom_im[469] = -9'd125;
    assign  twf_rom_re[470] = -9'd40;   assign  twf_rom_im[470] = -9'd122;
    assign  twf_rom_re[471] = -9'd50;   assign  twf_rom_im[471] = -9'd118;
    assign  twf_rom_re[472] = -9'd60;   assign  twf_rom_im[472] = -9'd113;
    assign  twf_rom_re[473] = -9'd70;   assign  twf_rom_im[473] = -9'd107;
    assign  twf_rom_re[474] = -9'd79;   assign  twf_rom_im[474] = -9'd101;
    assign  twf_rom_re[475] = -9'd87;   assign  twf_rom_im[475] = -9'd94;
    assign  twf_rom_re[476] = -9'd95;   assign  twf_rom_im[476] = -9'd86;
    assign  twf_rom_re[477] = -9'd102;  assign  twf_rom_im[477] = -9'd78;
    assign  twf_rom_re[478] = -9'd108;  assign  twf_rom_im[478] = -9'd68;
    assign  twf_rom_re[479] = -9'd114;  assign  twf_rom_im[479] = -9'd59;
    assign  twf_rom_re[480] = -9'd118;  assign  twf_rom_im[480] = -9'd49;
    assign  twf_rom_re[481] = -9'd122;  assign  twf_rom_im[481] = -9'd39;
    assign  twf_rom_re[482] = -9'd125;  assign  twf_rom_im[482] = -9'd28;
    assign  twf_rom_re[483] = -9'd127;  assign  twf_rom_im[483] = -9'd17;
    assign  twf_rom_re[484] = -9'd128;  assign  twf_rom_im[484] = -9'd6;
    assign  twf_rom_re[485] = -9'd128;  assign  twf_rom_im[485] = 9'd5;
    assign  twf_rom_re[486] = -9'd127;  assign  twf_rom_im[486] = 9'd16;
    assign  twf_rom_re[487] = -9'd125;  assign  twf_rom_im[487] = 9'd27;
    assign  twf_rom_re[488] = -9'd122;  assign  twf_rom_im[488] = 9'd37;
    assign  twf_rom_re[489] = -9'd119;  assign  twf_rom_im[489] = 9'd48;
    assign  twf_rom_re[490] = -9'd114;  assign  twf_rom_im[490] = 9'd58;
    assign  twf_rom_re[491] = -9'd109;  assign  twf_rom_im[491] = 9'd67;
    assign  twf_rom_re[492] = -9'd103;  assign  twf_rom_im[492] = 9'd76;
    assign  twf_rom_re[493] = -9'd96;   assign  twf_rom_im[493] = 9'd85;
    assign  twf_rom_re[494] = -9'd88;   assign  twf_rom_im[494] = 9'd93;
    assign  twf_rom_re[495] = -9'd80;   assign  twf_rom_im[495] = 9'd100;
    assign  twf_rom_re[496] = -9'd71;   assign  twf_rom_im[496] = 9'd106;
    assign  twf_rom_re[497] = -9'd62;   assign  twf_rom_im[497] = 9'd112;
    assign  twf_rom_re[498] = -9'd52;   assign  twf_rom_im[498] = 9'd117;
    assign  twf_rom_re[499] = -9'd42;   assign  twf_rom_im[499] = 9'd121;
    assign  twf_rom_re[500] = -9'd31;   assign  twf_rom_im[500] = 9'd124;
    assign  twf_rom_re[501] = -9'd20;   assign  twf_rom_im[501] = 9'd126;
    assign  twf_rom_re[502] = -9'd9;    assign  twf_rom_im[502] = 9'd128;
    assign  twf_rom_re[503] = 9'd2;     assign  twf_rom_im[503] = 9'd128;
    assign  twf_rom_re[504] = 9'd13;    assign  twf_rom_im[504] = 9'd127;
    assign  twf_rom_re[505] = 9'd23;    assign  twf_rom_im[505] = 9'd126;
    assign  twf_rom_re[506] = 9'd34;    assign  twf_rom_im[506] = 9'd123;
    assign  twf_rom_re[507] = 9'd45;    assign  twf_rom_im[507] = 9'd120;
    assign  twf_rom_re[508] = 9'd55;    assign  twf_rom_im[508] = 9'd116;
    assign  twf_rom_re[509] = 9'd64;    assign  twf_rom_im[509] = 9'd111;
    assign  twf_rom_re[510] = 9'd74;    assign  twf_rom_im[510] = 9'd105;
    assign  twf_rom_re[511] = 9'd82;    assign  twf_rom_im[511] = 9'd98;


endmodule
